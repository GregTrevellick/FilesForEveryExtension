Foo bar CKT