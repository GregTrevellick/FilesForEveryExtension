Foo bar BSV