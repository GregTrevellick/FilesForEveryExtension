Foo bar VHD