Foo bar CDL