Foo bar SVH