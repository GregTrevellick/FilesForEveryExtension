Foo bar LEF